library verilog;
use verilog.vl_types.all;
entity bancoRegistradores_vlg_vec_tst is
end bancoRegistradores_vlg_vec_tst;
